netcdf test {

 dimensions:
   n = 10, time = unlimited;

 variables:
   int n(n);
   int time(time);
   real var(time, n);

 data:
   time=1;
   n=11,12,13,14,15,16,17,18,19,20;
   var=1.1,1.2,1.3,1.4,1.5,1.6,1.7,1.8,1.9,2.0;
}
